module main

const version = '1.1.0'
