module common

pub struct Empty {}
