module main

const version = '1.4.0'
