module main

const version = '1.0.1'
