module main

const version = '1.3.2'
