module main

const version = '0.1.0'
