module main

const version = '1.2.0'
