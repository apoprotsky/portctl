module main

const version = '1.5.0'
